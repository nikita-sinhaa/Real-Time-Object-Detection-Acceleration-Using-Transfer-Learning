-- Placeholder testbench for bbox_filter.vhd
